//
// wshb2avl.sv
// @brief : 
//     A wishbone to avalon bridge
//     The avalon interface uses only burst mode for both read and write
//     For Read requests, we use a fifo to store the entire readdata burst 
//     since the avalon readdata has to be consumed as soon as the readdatavalid is asserted.
//
//     Using burst mode for write was required since we noticed an abnormal behaviaral of the DDR3 
//     simulation model when a  sequence of write requests occur with no burst mode.
//     The DDr3 simulation model was generated by qsys soc_system testbench generation.
//
`default_nettype none
module wshb2avl 
#(
    parameter ADDR_WIDTH   = 32,
    parameter DATA_WIDTH   = 32,
    parameter AVL_BURST_LENGTH = 8
)
(
    wshb_if.slave wshb_ifs,
    avl_if.master avl_ifm,

//--- Just for Debug
//   output wire w2a_rsp_fifo_full,
//   output wire w2a_rsp_fifo_empty,
//
//   output wire w2a_wr_fifo_full,
//   output wire w2a_wr_fifo_empty,
//
//   output wire w2a_avl_write,
//
//   output wire fsm_wb_id,
//   output wire fsm_wb_write,
//   output wire fsm_wb_read,
//   output wire fsm_wb_flush,
//
//   output wire fsm_avl_id,
//   output wire fsm_avl_read,
//   output wire fsm_avl_write,
//
//--- 
    input wire [31:0] img_addr
);

wire  [ADDR_WIDTH+DATA_WIDTH-1:0] wr_fifo_rdata;
wire  [ADDR_WIDTH+DATA_WIDTH-1:0] wr_fifo_wdata;
logic wr_fifo_write;
wire  wr_fifo_read;
wire  wr_fifo_full;
wire  wr_fifo_alfull;
wire  wr_fifo_empty;
wire  wr_fifo_alempty;

wire  [ADDR_WIDTH+DATA_WIDTH-1:0] read_fifo_rdata;
wire  [ADDR_WIDTH+DATA_WIDTH-1:0] read_fifo_wdata;
logic read_fifo_write;
wire  read_fifo_read;
wire  read_fifo_full;
wire  read_fifo_alfull;
wire  read_fifo_empty;
wire  read_fifo_alempty;

wire valid_read_req  = wshb_ifs.cyc && wshb_ifs.stb && !wshb_ifs.we;
wire valid_write_req = wshb_ifs.cyc && wshb_ifs.stb &&  wshb_ifs.we;

logic [ADDR_WIDTH-1:0] r_addr;
logic [ADDR_WIDTH-1:0] r_waddr;
// max burst = 256 beats
logic [7:0] r_burst_count;
logic [7:0] r_wburst_count;
logic [7:0] r_burst_avl_wr;

logic wb_write_set, avl_write_rst, wb_avail_write;
logic avl_read_set, wb_read_rst  , avl_avail_read;

// RS-flip-flop used as a communication buffer between wishbone and avalon fsms
// It is set by wishbone fsm to request avalon write
// it is reset by avalon fsm when write burst complete (burst_counter = 0)
sr_ff
sr_ff_wr
(
    .clk(wshb_ifs.clk),
    .reset(wshb_ifs.rst),
    .set(wb_write_set),
    .rst(avl_write_rst),
    .state(wb_avail_write)
);

// RS-flip-flop used as a communication buffer between avalon and wishbone fsms
// it is set by avalon fsm when first read data available
// It is reset by wishbone fsm when read burst complete (read fifo empty)
sr_ff
sr_ff_rd
(
    .clk(wshb_ifs.clk),
    .reset(wshb_ifs.rst),
    .set(avl_read_set),
    .rst(wb_read_rst),
    .state(avl_avail_read)
);
//---- Avalon
typedef enum logic [1:0] {AVL_IDLE, RD_BURST, WR_BURST} avl_fsm;
avl_fsm r_avl_state;

wire match_write_addr = wshb_ifs.adr == r_waddr;

assign avl_write_rst = (r_avl_state == WR_BURST) && !avl_ifm.waitrequest && (r_burst_count == '0);
assign avl_read_set = (r_avl_state == RD_BURST) && avl_ifm.readdatavalid && (r_burst_count == AVL_BURST_LENGTH - 1);

always_ff @(posedge wshb_ifs.clk)
    if(wshb_ifs.rst) 
    begin
        r_avl_state   <= AVL_IDLE;
        r_addr        <= '0;
        r_burst_count <= '0;
    end
    else
        case (r_avl_state)
            AVL_IDLE:
                if(wb_avail_write)
                begin
                    r_burst_count <= r_burst_avl_wr - 1'b1;
                    r_avl_state   <= WR_BURST;
                end
                else if(valid_read_req && !avl_ifm.waitrequest && !avl_avail_read)
                begin
                    // send avl read request
                    r_addr        <= wshb_ifs.adr;
                    r_burst_count <= '0;
                    r_avl_state   <= RD_BURST;
                end

            WR_BURST:
                if(!avl_ifm.waitrequest)
                begin
                    if(!wr_fifo_empty)
                    begin
                        // wr_fifo_read = 1
                        if(r_burst_count == '0)
                            r_avl_state <= AVL_IDLE;
                        else
                        begin
                            r_burst_count <= r_burst_count - 1'b1;
                        end
                    end
                end

            RD_BURST:
                if(avl_ifm.readdatavalid) 
                begin
                    // write fifo (readdata, r_addr)
                    if(r_burst_count == AVL_BURST_LENGTH - 1) // &&
                        r_avl_state <= AVL_IDLE;
                        // avl_read_set = 1
                    else
                    begin
                        r_addr        <= r_addr + 4'h4;
                        r_burst_count <= r_burst_count + 1'b1;
                    end
                end

            default:
                r_avl_state <= AVL_IDLE;
        endcase

assign read_fifo_write  = (r_avl_state == RD_BURST) && avl_ifm.readdatavalid;
assign read_fifo_wdata  = {r_addr, avl_ifm.readdata};

assign wr_fifo_read       = (r_avl_state == WR_BURST) && !avl_ifm.waitrequest;

assign avl_ifm.address    = img_addr + ((r_avl_state == WR_BURST) ? wr_fifo_rdata[ADDR_WIDTH+DATA_WIDTH-1:DATA_WIDTH] : wshb_ifs.adr);
assign avl_ifm.read       = (r_avl_state == AVL_IDLE) && !wb_avail_write && valid_read_req && !avl_avail_read;
assign avl_ifm.write      = (r_avl_state == WR_BURST) && !wr_fifo_empty;
assign avl_ifm.writedata  = wr_fifo_rdata[DATA_WIDTH-1:0];
assign avl_ifm.byteenable = '1;
assign avl_ifm.burstcount = (r_avl_state == WR_BURST) ? r_burst_avl_wr : AVL_BURST_LENGTH;

//---- wishbone 
typedef enum logic [1:0] {WB_IDLE, WB_FIFO_WRITE, WB_FIFO_READ, WB_FIFO_FLUSH} wb_fsm;
wb_fsm r_wb_state;

wire match_read_addr = wshb_ifs.adr == read_fifo_rdata[ADDR_WIDTH+DATA_WIDTH-1:DATA_WIDTH];

always_ff @(posedge wshb_ifs.clk)
    if(wshb_ifs.rst)
    begin
        r_wb_state     <= WB_IDLE;
        r_waddr        <= '0;
        r_wburst_count <= '0;
        r_burst_avl_wr <= '0;
    end
    else
        case (r_wb_state)
            WB_IDLE:
                if(valid_write_req)
                begin
                    r_waddr        <= wshb_ifs.adr;
                    r_wburst_count <= '0;
                 // r_burst_avl_wr <= '0;
                    r_wb_state     <= WB_FIFO_WRITE;
                end
                else if(valid_read_req) 
                    r_wb_state <= WB_FIFO_READ;

            WB_FIFO_WRITE:
                if(!wr_fifo_full)
                begin
                    if (valid_write_req && match_write_addr)
                    begin
                        // fifo_write = 1
                        r_waddr        <= r_waddr + 4'h4;
                        r_wburst_count <= r_wburst_count + 1'b1;
                    end
                 // else if ((valid_write_req && !match_write_addr) || valid_read_req)
                    else if (valid_write_req && !match_write_addr)
                         begin
                             if(!wb_avail_write)
                             begin
                                 r_burst_avl_wr <= r_wburst_count;
                                 r_wb_state     <= WB_IDLE;
                             end
                         end
                end
                else if(!wb_avail_write) // wr_fifo_full
                begin
                     r_burst_avl_wr <= r_wburst_count;
                     r_wb_state     <= WB_IDLE;
                end

            WB_FIFO_READ:
            if(avl_avail_read)
            begin
                    if(read_fifo_empty)
                    begin
                        // avl_read_reset = 1
                        r_wb_state <= WB_IDLE;
                    end
                    else if ((valid_read_req && !match_read_addr) || valid_write_req)
                            r_wb_state <= WB_FIFO_FLUSH;
            end

            WB_FIFO_FLUSH:
                if(read_fifo_empty) 
                    // avl_read_reset = 1
                    r_wb_state <= WB_IDLE;
                    // read fifo until empty
            default:
                r_wb_state <= WB_IDLE;
        endcase

 logic wb_read_ack;
 logic wb_write_ack;

// assign wb_write_set = (r_wb_state == WB_FIFO_WRITE) && (wr_fifo_full || (valid_write_req && !match_write_addr) || valid_read_req);
 assign wb_write_set = (r_wb_state == WB_FIFO_WRITE) && (wr_fifo_full || (valid_write_req && !match_write_addr));
 assign wb_read_rst  = ((r_wb_state == WB_FIFO_READ) && avl_avail_read && read_fifo_empty) || (r_wb_state == WB_FIFO_FLUSH);

 assign wr_fifo_write = (r_wb_state == WB_FIFO_WRITE) && valid_write_req && match_write_addr;
 assign wr_fifo_wdata = {wshb_ifs.adr, wshb_ifs.dat_ms};

 assign wb_write_ack  = (r_wb_state == WB_FIFO_WRITE) && valid_write_req && match_write_addr && !wr_fifo_full;

 assign read_fifo_read = (r_wb_state == WB_FIFO_READ) && avl_avail_read && valid_read_req && match_read_addr; 
 assign wb_read_ack   = read_fifo_read && !read_fifo_empty;

 assign wshb_ifs.ack = wb_read_ack || wb_write_ack;
 assign wshb_ifs.dat_sm = read_fifo_rdata[DATA_WIDTH-1:0];
 assign wshb_ifs.err = 1'b0;
 assign wshb_ifs.rty = 1'b0;

wire read_fifo_rst = wshb_ifs.rst || (r_wb_state == WB_FIFO_FLUSH);

sync_fifo
#(
    .WIDTH(ADDR_WIDTH+DATA_WIDTH),
    .DEPTH(8)
)
wr_fifo_i
(
    .clk(wshb_ifs.clk),
    .reset(wshb_ifs.rst),
    .write(wr_fifo_write),
    .wdata(wr_fifo_wdata),
    .read(wr_fifo_read ),
    .rdata(wr_fifo_rdata),
    .empty(wr_fifo_empty),
    .full (wr_fifo_full),
    .almost_full (wr_fifo_alfull),
    .almost_empty(wr_fifo_alempty)
);

sync_fifo
#(
    .WIDTH(ADDR_WIDTH+DATA_WIDTH),
    .DEPTH(AVL_BURST_LENGTH)
)
read_fifo_i
(
    .clk(wshb_ifs.clk),
    .reset(read_fifo_rst),
    .write(read_fifo_write),
    .wdata(read_fifo_wdata),
    .read(read_fifo_read ),
    .rdata(read_fifo_rdata),
    .empty(read_fifo_empty),
    .full (read_fifo_full),
    .almost_full (read_fifo_alfull),
    .almost_empty(read_fifo_alempty)
);

//--- Just for Debug
// assign w2a_rsp_fifo_full  = read_fifo_full;
// assign w2a_rsp_fifo_empty = read_fifo_empty;
// assign w2a_wr_fifo_full   = wr_fifo_full;
// assign w2a_wr_fifo_empty  = wr_fifo_empty;
// assign w2a_avl_write      = wb_avail_write;
//
// assign fsm_wb_id    = (r_wb_state == WB_IDLE);
// assign fsm_wb_write = (r_wb_state == WB_FIFO_WRITE);
// assign fsm_wb_read  = (r_wb_state == WB_FIFO_READ);
// assign fsm_wb_flush = (r_wb_state == WB_FIFO_FLUSH);
//
// assign fsm_avl_id    = (r_avl_state == AVL_IDLE);
// assign fsm_avl_read  = (r_avl_state == RD_BURST);
// assign fsm_avl_write = (r_avl_state == WR_BURST);
//--- 

endmodule


